library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;  
entity Instruction_Memory is
	port (
		Read_Addr: in std_logic_vector(31 downto 0);
		Instr : out  std_logic_vector(31 downto 0)
	);
end Instruction_Memory;

architecture Behavioral of Instruction_Memory is
type ROM_type is array (0 to 31) of std_logic_vector(31 downto 0);
constant rom_data: ROM_type:=(
		"10101100000000000000000000000000",--SW $0,0($zero)  $s0=5 donc #5 <= 5 
		
		"10001100000011100000000000000000",--LW $14,0($zero)	$14 <= #5=5
		
		"00100001110011100000000000000010",--Addi $14,$14,2  $14=5+2=7 
		
		
      "00000000111010000011000000100000",--Add  $6,$7,$8    $6 = 7+ 8 =15
		"00000000110001010001100000100000",--Add  $3,$6,$5    $3 =15+ 5 =20
		"00000000001001100000000000100000",--add  $0,$1,$6 	$0 = 1+15 =16
		
		"00000000000000000000000000000000",
		
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		
		
		--"10001100000011100000000000000000",--LW $14,0($zero)	$16=#16=16   Change $16 here to smtg else
		
		--"11111100000000000000000000000000",--NOP
		
		--"00100001110011100000000000000010",--Addi $14,$14,2  $14=16+2=18 
		
		--"00100001110011100000000000000010",--Addi $16,$16,2  $14=16+2=20
		
	--	"00100001110011100000000000000010",--Addi $16,$16,2  $14=16+2=22 
		
		--"00100001110011100000000000000010",--Addi $16,$16,2  $14=16+2=24 
		
		--"00100001110011100000000000000010",--Addi $16,$16,2  $14=16+2=26 
		

		
		
		--"00000000000000000000000000000000",--NOP	
	   --"00000000000000000000000000000000",--NOP
	   --"00000000000000000000000000000000",--NOP	
		
		--"00100010000100000000000000000010",--Addi $16,$16,2  $16=8+2=10 
		
		--"00000000111010000011000000100000",--Add  $6,$7,$8 =15
		
		--"00000000110001010001100000100000",--Add  $3,$6,$5 =15+5=20
		
		"00000000001000100000000000100000",--add $0,$1,$2=3 
		
		"00100010000100000000000000000010",--Addi $16,$16,2  $16=8+2=10
		
		"00000001010010110100100000100000",--add $9,$10,$11=21
		
		"00000000111010000011000000100000",--Add  $6,$7,$8 =15
		
		--"00000000110001010001100000100000",--Add  $3,$6,$5 =15+5=20
		
		--"00000000001000100000000000100000",--add $0,$1,$2=3 
		
		--"00100010000100000000000000000001",--Addi $16,$16,1   10+1=11 

		--"00000000000000000000000000000000",
		
		--"00000000000000000000000000000000",
		
		--"00000000000000000000000000000000",
	
		--"00000000000000000000000000000000",
		
		--"00000010000010011000000000100000",--Add  $s0,$t1,4
		--"10101100000010000000000000000000",--SW $t0,0($zero)
		
		
		--"00000000000000000000000000000000",
		
		--"00000000000000000000000000000000",
		
		
		--"10001100000100000000000000000000",--LW $s0,0($zero)
		
		
--		"00100010000100000000000000000000",--Addi $s0,$s0,0
--		
--		"00100001001010010000000000000100",--Addi $t1,$t1,4
--		
--		"00100001000010000000000000000011",--Addi $t0,$t0,3 
--		
--		"00000010000010001000000000100100",--And  $s0,$s0,t0
--		"00010001000100000000000000000010",--beq  $t0,$s0,+2 -3(1111111111111100)
--		"00000010000010011000000000100010",--sub  $s0,$t1,4	
--		"00001000000000000000000000000010",--j    2
--		
--			
--		"00000010000010011000000000100010",--sub  $s0,$t1,4	
--		"00000010000010011000000000100010",--sub  $s0,$t1,4	
		--"00000000000000000000000000000000",
		--"00000000000000000000000000000000",
		--"00000000000000000000000000000000",
		--"00000000000000000000000000000000",
		--"00000000000000000000000000000000",
			
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
	
	
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000"
  );

begin
	Instr <= rom_data(to_integer(unsigned(Read_Addr)));
end Behavioral;


















--library IEEE;
--use IEEE.STD_LOGIC_1164.ALL;
--USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--
--entity Instruction_Memory is
--
--	PORT (address: in STD_LOGIC_VECTOR(31 DOWNTO 0);
--	
--			data: out STD_LOGIC_VECTOR(31 DOWNTO 0));
--			
--end Instruction_Memory;
--
--architecture Behavioral of Instruction_Memory is
--
--TYPE rom IS ARRAY (0 TO 256) OF STD_LOGIC_VECTOR(31 DOWNTO 0);  -- 1kbytes of memory
--
--	CONSTANT imem: rom:=(
--   "1000000110000000",
--   "0010110010001011",
--   "1100010000000011",
--   "0001000111000000",
--   "1110110110000001",
--   "1100000001111011",
--   "0000000000000000",
--   "0000000000000000",
--   "0000000000000000",
--   "0000000000000000",
--   "0000000000000000",
--   "0000000000000000",
--   "0000000000000000",
--   "0000000000000000",
--   "0000000000000000",
--   "0000000000000000"
--  );
--
--	
--	begin
--	
--	data<=imem(TO_INTEGER(address));
--	
--end Behavioral;