-- An array of instruction 32*32, the output is the instruction at the read address index.

library IEEE; use IEEE.STD_LOGIC_1164.ALL; USE IEEE.numeric_std.all;  
entity Instruction_Memory is
	port (
		Read_Addr: in std_logic_vector(31 downto 0);
		Instr : out  std_logic_vector(31 downto 0)
	);
end entity;

architecture arch of Instruction_Memory is

type ROM_type is array (0 to 31) of std_logic_vector(31 downto 0);

constant rom_data: ROM_type:=(

		"00000001101101010100000000100000",  --add $t0,$t5,$s5
		"00000001101101010100000000100010",  --sub$t0,$t5,$s6
		"00000001101101010100000000100100",  --and$t0,$t5,$s7
		
		"00000001101101010100000000100000",
		"00000001101101010100000000100010",
		"00000001101101010100000000100100",
		
		"00000001101101010100000000100000",
		"00000001101101010100000000100010",
		"00000001101101010100000000100100",
		
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000"
  );

begin
	Instr <= rom_data(to_integer(unsigned(Read_Addr)));
end arch;

--
--		"00100001000010000000000000000011",--Addi $t0,$t0,3  // t0=8+3=11
--		
--		"10101101000010000000000000000000",--SW $t0,0($t0)
--				
--		"10001101000100000000000000000000",--LW $s0,0($t0)  // s0=11
--
--		"00000010000010011000000000100000",--Add $s0,$s0,$t1  // s0=11+9=20
--
--		"00000011101010111000100000100010",--sub $s1,$r29,$t3  //s1= 29 - 11 = 18	//s1 = 29 - 9 = 20		
--
--		"00010010001100000000000000000010",--beq  $s1,$s0,+2 //18!=20 => no branch  //20==20 => branch taken, program counter goes to nop instructions.
--
--		"00000001011010010101100000100100",--And  $t3,$t3,t1 // t3 = 11 and 9 = 9
--
--		"00001000000000000000000000000100",--j    4